`ifdef RTL
	`define CYCLE_TIME_clk1 17.1
	`define CYCLE_TIME_clk2 10.1
`endif
`ifdef GATE
	`define CYCLE_TIME_clk1 47.1
	`define CYCLE_TIME_clk2 10.1
`endif


module PATTERN
`protected
c\SMOd9UD>H-CeBgL-M5&53P9JJQ3I7@&=K?TXI;_CR6=Q6?Y.K(-),NO#02?-<=
^[9:IJ8#Mg+)5Y\ZBR0KHWYQU#@YI7beB8)VB(SLJgbV4Q@5]c.E,U08)Q:M9=FX
L:<SbWcbRaeX_-dG/T(X@/c(bN;LP.(cgHZ\(4#G51f7V:@)I4A0/E@T(f)ABBV,
Cc(C<dbe5<?OKVU]QQc7;9_ZfX&K3[cJfR(:fFD&^-8/:XKE..ORf;.B,/TEC?^U
I#H9&N#@<:E.WWd35T)X6\&1Ve7<9D>]gL7YTBC9+.;21.@.aS7:K=A/)c[&OUF(
2(=O7TKeV/:9/WUXffVRSGTU@:4;L-:<89^De0E0Y9JA/[RD5Eg5WFA&;R[C^61S
1HcRCDSWIHBK3[VF&][]2Xg3(Fd#5G[#-L(SA-0J@6B3L^\^A.2XV940+0EC?,GA
M>0CYUeb#X=[Me_]658L@V10&/gSQbJcN>eYA.\NA6;-:XTVXHfbXg+#;PRL]8)F
AV8HX.=F=8AX6AOP:>aTH[G3J2:I06]>).F0_3A/b:-&Jb4PCPHDQJge+fc7-\EV
+A;:7>)[76S^O(@TX+HUXgWD-?4gGfUOIcbEF9K,BGG<=g8>1QUQGcU@R_6\NF,e
7,1/7aA]AQdQ1YS0E5E_fBMP)c8(XUCTR\7ISFQ@]&EfgUgV+8NI(OcQ>B978YLY
C5G:W0H=T8K\-_g]:2\;F-AFfeT[ce0.^R1F6B+N<1@KE2\SdY<1YTA6P(8./9cQ
9R#,0-fa7#eFM5R@,AOY\YJND4dB=.5cWF.I;3^T)#IZ(WX:ALdVHAW0&4^/.+b:
f#cVDO83WL\W(35T,,WTM?c+;A\G)S+5Ib)E](SXY780,-0_VG5a8[eD)d\B8QUC
AfE3?<W<T8R5\(P/M0=6R?H?M25/T<^RgK/=g8RU]X60&?ON3=f)DM8XL0<;FWR(
.>)@=76-;aZ1(2C9,QW#f86>McUPgBG\E;>NMd)JTH=/fgb-ea+4MR:aD#VMH2OJ
\J>-6#_F7dM1>ITS5caFT4[8F5+f\>\\41JJP86:b83(N([#Q<]aU:b5Q>=8VP7J
Sa,-d^-;G\JFRGYR4=UY[5-@JT:E;W-:?M()3;Af<D]_[_T(61,IGFLPM8><dGMg
-VIK&@GcV_DGSIR;Y<J7Wc/PM@6Y21VDbUZI::7@NOE<JV@DXc@RR6W?NX4?1^0S
#>9B9/@Q@3e<A??_1@35_cO4X;RaH4(8EXL<caCS+e5<J:Y^cEg[OG>@.AFL03XW
7JgP-/>WJG2_O[B9bAG>YJ^gV0G;:GX7MF4RYfE-S@f9?69(AC@WOb8;+ROJ;3/(
,eG8A;E@UcE[S,&3e/QZQZ^17=dfW-FZ=YY1>((@HgcMMAcbVf)3\<@/7M:7-f@<
6a?gYUG9I.AOY+C]L]RJ5I(CA?K(VK@f@<8+G53?K-ZQH\LSG_;/eIcJCT1PI1EG
#3cQNUN[EGWW#T0P#LOXJ?@VR,-O\NUKS):28XD27a)Ee^+30a?^(Yd+@=g+[VM0
e[EWZ_cZT8g2]2bTOC^]bdJ-)_J@V)/de;R[]:JR_0IL[)B3@L.QD<4^(8@[]Z&]
S(A3PSNAD<M_^I0^RQSU_gg#6WZN[;R&aT.b4EH0UJWg3YR,>4KJM?J]Gdfd?XK5
:g,?,-d.TU[RJ2+&cC1eL0EL<QV_-4OMba==P]]]7dII&AK],7/N,K/KZK+K->[G
L9X^]1JYG]3))Me#A&6NeISV[>F\[:WE@<+b-ZOGWZ=cGC4<^e,2UNJWHV3TKV/C
CY_)TE5E7eC^5Fe5dAbJ>:DUJ[)8PE+g7\L8H2PWWA7\G-&=KaPO@OYEV^A;g>@;
YX;Y9](_>f1N1b_Le7SJeRC6Ac5d8JC3P,We==GcR=4ZWS>XO->]KPbDAW?-M@+K
\VNa@9O?NaZ[^a10G7,c&^01?,IF8;IbK(6V0gQ2eK5<6=^&P2@C42d#:0#.aTd<
c,:V[W<c757bbWXCO0#dC+(6bJDL4R>BZS+W05A[@cb(&3Jd^G?:8_RXU7_6NT[T
WB70[28TQYd\X41#(/SW(04QV:]TdM:&4U2W-fN)SXNG4DLYg83(AZH6]Z^_Y&?4
cQY_8_D&9&YZ#(BDN2]W2W2^cU5dMV6U7aQH>;52f;+/?(6Cc)R^I1178.FS9XAG
g_P<CPbL,FK?L,_/Z#P5gMYb;,7MWN5AHXJ.O@1#;OC)Z_,#NgQfb)Uf6CNJ3g^<
d>T4VaUHH+8Mb-,U@HN/G\a==4ecO90(QQ[.&edVI:6J?e<2]5C8L,:U2#^EOEd[
)d8SGNLJQDF>DW?Y#R@N?&cda5GZ&#++J=S8Z00bOaP#;]Td3QgZdf[O;:JK)RgR
Q(T1<M5ad_dFbK,A>9+VeeQOg3P^d[EP?:Z?7^NV@MJ0X)H4e#/\IfgeKGO,11M)
0faUJCX7Y+BI+M97G@C9g^[-:gWcDZHa^23MDST51ZQKW;=e6+TcfM5[1@9EH(]K
,SXO(VRg3U[OD)WI?df6UTZ#9RQ6M.4IEZ)La7JDIF?\,]6:cX)-8F5YQ:XZZ<FV
E+9gObB8W)/>f(7FO+5#[?I2;-EB]4_M:b9[dF,O.DG6eF4.+@SeV;#5a3B1N5)^
(]9JB]fIX8O5.TecT7eB+gP[=Ia4LUB5,\NS_GM6>5318:IMF;dXZ<M(72:+c/MZ
S#RWTTI@5BA)ETD#;a)^^E+JcN@8JJGK9;^;cNNB2X.DgWY/.F+30=1c\IX)cEe@
[\BL.,A\4V5c8-bSaIUb@84791CDMRMfZ[VU[M,bJ:NO_G89O(^\Xd=949\^#7,;
2c[3J2fQG71E^(?dOBB4,1AP8IQ.41;OOQ2f25HP-.+;KHOb14c(Y-5Q]>EPKI50
Z37L&b?2W@[(-@_L(R(-aA4Yc+9^A0=4He7A:(1_R=E2@E#<W<[I4M=?c]@#bXL(
M.V/f=R&cH6dHA#a4SHObDDWF>Y2KFKHNId_+XaJ,?Ia01X5^-><c<<-V-bM8Zff
0SV:Z]=64SOL=),IU75FK9XA#T-b/RII&(],#F0@:3B:]O11B<O0b2KMRL+;?YFg
J.@,VU.\4]Ud7-XbDfD3OBI&Feb(dW2eHU027(GXfV[Y_I+7?a,1K.E0RU(>X1BB
VaPc7]<[aO3ZSSW)VabL56/gEC>dg7eAa8D#U]GVb0I\H<9JRM?MCL_J4C<>IaXf
79Ra(a8B-0E&;/c:OEDcTf#NY\c)PT<-b32XEQF<562]gI<.W]ITD&1J_51C?0I0
3Gb,1,\4TYNJbK,bU-,a(_JC0^PG=BNL).GeZ36R.-]G+#48U1CMF7&SR-(JI.6D
)SgZ>dXA()M077a.)g9D2S]>fc@Se^9F64_Z<>Hb0:&7EY2SL7:6560>0&F?PCD1
6=PeFIPBXCL85V<8=dK_S62KB43\).S(GUEADeFg),1OA;ab1Ffbf)D?2IgfZe:-
,2P:b>XW?FAeN^CY>1f4VVT4D#RQL^/MD.bOe76&)X@@:@E0UaX<OZQgC<4Pd9?F
YPS//.Hd5RV+.LB<M=T=D&ec\JN0_#SKFc(8K=6IH4MM_Y>F\bRNH;YTaNdY)KA.
YH9NV4U7DWbH6TTIHS?2aeLc;GS[T5\&S>Af&[E)Q#JCbE<>IDWL/:I\7F)R-V^;
eW6,?COPBD6OSR@Of&D&-M=GbM5::CVF610d03V_g\Mg<_BWKR1F-5I@6&+(,FS&
=1\U=c_=92e]0]c?a6CWbeecd=Zd,1WM;Z\?S=L/-=AG#2Sc^I4S\:@=Y,6X3_._
K;=R<J5-Ia[\_K<2W,&24Y<.Z6)KJ:9N;>YD8cfSaL3V9LL?bSeCg1RM3DDR/=EI
A,]SRQ]d#RXb<AL^c+NQ6CXM0IDGQ=18f(7\0g<<+Kg\&ZeU1U8VU8/.&)cQ-A;[
GJ>dfQ+MaIcG?/ee-CY=<X:3U)cA4&9^NWU3fFNS6cCR_PUB+Y3O9Eb^;P==CVNJ
L1]e2(^+AX0.TK20,(ALHCb1/;+20:R4#3b/3U83.)CgM>I:G2[]3f>N=5XEF7/K
^:BbYb7<Q35B)IB:cfV3Y3;b0<?YPCa,M^4_5]1N>YH@]=2@#cUHKY4TB_/=g<X8
//cP#(;4f1f.7J3/8:Q[:#,>O\^GLJ.5_ggbQ0P^MGM5dMWFGQ5/CRT71UNYd(GM
>:V/aW[.OH?F=NRHDLb?6>,US\R[@?(WR8(g14E[&WVg8Y#^MA]dX=3N0P,D&..(
ITV\M896B7XJQP2c_HKX4IYH:f.aa#XEW[3aI/?;MS_J&K&_#SCBIBH:#[g>gf02
]Xd;]S,(JGc8_I&C_Mf3B95WP\g/.MC6IS12&0U.YWKZHPI))fe,5DBUU?-IX+.>
QD,S-V@AV-9J2[Hd)QFFK(-a/.IeLbJ1ZLg&<=2+#ZTIE3b#g>55[5cI9?]HAIf,
2BP4#MSCDG\J)CX_C[WRT#F5+L96LCTLZPg>-_86\6Mg=/E8Z=,94N;A9G<c)b6g
-LUTeQ:WJV52Jbc;]G3-L3T9;^T-W^3H6/6Tga<[>eD4?,<NY41LURJNR)-K>1#A
);Mdb;<U#AXZ1,_HA_TOAgH1eH@I/b?&;gKPT+1>-;7]H]X9I:e)a@I1DYP>N@^Y
IJd50L/-a4G:NgC:C5ZJO0LXeEc-UgZI5b@ZW)cM:;f0AW#BCC(#A1</.I8E?\/;
5f5)JYZA-6#J38?O#.@,CGJ4.-/bQDXT3_@c2UO,4H<N;MY2-a#_(1BKO8T7@Q<+
XDTdB/ab.+K(G;Tf3PDI5<]]&Z-48-YJ\<@f/08fQQ^TEBM3.#WaH\0,)4;]4J\+
.U&9?CPf.G:4(0K<-5+-J,g?0bM1(CN^]<2P/,_>V7_>DLI_TYXKFg#F)@I#_Lf@
3[QeJ3,^ca<V7CB.IWPFcI_S8C2?D>b4>9/TY-]((113eKCX5.,?cD:K?JT<MCJ>
;VXaCMd+@HVB?^CYUQ#/Ta>,6.TC+@IBW\8SGAXU?4VET:ZM48Va_]FJ]\S0QB3T
gO:8PF_af;+K;BH.e?KK^+J@0cJB#]HQ5N-#U:.D3IZ0b>(EXXWIAg<8_QC&EWY>
Z18M[4eLOWP/1,fUTOO8@MWb^DbZ8[f(Pb00@=d]W/+)=@e;O_X7Le#H[[-4],fW
?#<QM)aC^93;5[-](.ED\R@XN0\:3=0^K74@X53I6^./D2fDW:Rg=<Te3.K#KR,;
FJg#G29Y46;F4_:cV8I0.,VG;Q?0P02^H>JRg;J_F+?.9TK&?7<:YAWXJe1X9G=f
5IE&&PCN(e=X3&\L.V?A(Yc+>a5dP-c_>d&_88K15c23&W?9HX5PIaX@3J?8?a3,
EFF[&f>_GP;Q,9T0V?K](/LBQ=#V,#Y>f0a^100+(2I+,F55;MIYb+a&;35<dNT#
(E#GCX7N>f@MA_=C/I31?f_U;Q9?)6DL2,C5X?a7?TQcG07[19c>e/PA;\ROEI,E
@//&72OdOIDGFTC(IXS]?&?I^:[JaQ#IY];[.,T\:NPUb,^:85Zb7+JB)OG1a[5&
.U5O1b5RV1->5SdAS&/aJd9T/OGe;O;GP.]7B9[BG8Ab^B)3_6TD::K2@1^&/UYe
ec+?2FFK;L&W\TY<I;)a6:@S;?@a&_]L5X1E<OUaUH(3/-ad/CGAA1G][f#T:e>c
[K?67eg>:3D3eEVbDURg&^F>e#I\(OU?FSe-JGWFcANO&4JU9K>7PN((5?KX@QIF
^^DIbY=H6_S>TO=4.1B(\I\P8&CHc_1_-bG0K^HYC;[#GQg[8K/a1EfI990JS,:.
bZPK5A1T8TMYT\DXaIB#NaJ(B5XPK/R(e]a_APGEf,e::=_6M,A0X2c]BfgBWG1[
Z@:aM4:V-25=VI59HQ:22TC#ZWNBgd_;VN:E)[CZ3&dP?L,65\EV6CVaWe,IW87=
ff@SB]I52^Ee8\\EOM\ELX\1[QU>&OH9aD-[BL;gbBFZYOG)RQJGKY2ZM>FE.Z;J
aV[WbF9KRO:ae/W>F_9&:VYRDCN_G^QF;HU>,KG9[=5ZXf[A7;4,KCTBa.UQK-Y+
SYGVbK>f[@8[Na;LCb2R3>0Q8/BSOaB>VMOLHQOV[7X/LZ2KZ,SHVD;0Q7g?]IB,
/T&V)<Rc-aSR5&B5D7G5Pe>#ac_eb(/F..-26e?9(VZ7I^_.FSTU7LJ/,B]WN+TR
bU.OE?>W[cJ8(8L64DP)feER[I9gF^^\#\VZ84GDCTfM9(]^&]Y(I\[2+H7[b@N7
Y8)>DK;Kb&=PVe.#5T8_gg<YP<33[WUX/eGCNFa/JcLGVTAa<E)^ESfDBT<J]8gF
H7U._B4=5#ETBU:bRfFK&:\UN>F/&OHJG[Z_eU._>VL>J]XfP->3c:T;@3Lb7b/P
MRCK;^B6b2Z@;S.DNX.AO<dWRVA=>Gd(Z&U7Z8ZQ(LfKKWKQ/eTBP>ca[X1Ia0;[
6W^>UbBQ;QV\ZHJb76DAW^=HE/U#_3-8;?Y31X]X-.M3ASB2<dB^#.V4_S7<3a/(
Rd2J4NdbSJ+/5HFR8U1E9_M8cK+7,PO09,2EDc)87Z4,)2#CVbcb?g2.GD73G5f)
G?0W24FG2eb+]AD\,?&@ASF(0<Eb?1#Q73J]bOcHXUGA=a<;7/Yf_DIKg^4egT:P
.:5a#I(0a?eZZ4BV?^=6D_\5/]ML8-a40)36.Z1I<VTA?Z3/T\A6M#FW&7c(R2,8
[7XaYZ1O@-,W:KO0)5K1bJ4D03VQFEU7_f3HRc7dN,9AV>AQ\S?FfdLJc)OU>dXA
RJ/?WLY@U@8^TEfCU0]>(Y</6HaRE7]QVXAaO+UHFRG@3EO+<500[^]\BRRDS=bW
HK445?^UBEdR\0N)?Cc5K?>BB]HXGN..Y[ZJ4HfL=(d\,[;c8P@F=XDA2)a]QJ\I
b>\b@#Ugf2&G+_<_KD&gg(H@L;)/9J7A5EIUWc/<a\/:[9WJ&G2YSEb&_bJCF7.;
3J=Id_D9[.4L7Z>SRJLZb&1JTG9(,GYU39b(,?aRRdVA-.O#P8AJF<WG#31g=PK<
aIdN6E/>b5;[9+3gO/^>5WV8U\#g.I,W#,HCJGMRT.,V(7]J)&\X3XU+2</^?aZV
-9ccgTMVWdGWcQf1/@bLeLGg)Q@/62(5]KOeAFV>6AEUG8Na>c,UN9d#?9J?e_J+
K(4EC0]JF5YaLX0(NI+P-ER+a?dg,CS+2VZGSd^2<<g4-F:e\[V.H;gF0+/OJDW&
-GfeP9YPaRBgddS0;7MY1>^6/K<2>GIV8&A(I;6&TZf1Ca(DZ#1.MQFT->bCb\0=
M(bf2d_Q/IV/Kgf?eGQg^6fgHWGBJ+4>bP,O+\_[N:R;@d\Wa(<Tdg6>[<BZ<G.^
4M]7GCQ)-UJc&gV-H(8g(P_HdA#CJ(d4R<ZV(a(9e.:-O<52NBgI-d;^LK.bY;aO
#RC@L2>DFI?Z>E4:W8QAV=-6dPKDVTO0NOV<MW>:\_8KdWWBE#3^SVgFQLTX8#JT
Q9@5(R89B_;=\&0]0K).1Ga+5A5YK:[[SDgcO>>\OZL-;5X?EED_Y.M<&9;>1^ZO
\R.VK#[21dA^+XT+<ROYMT#;,Q^5afEB2?Ne6)RRJXE^KMg:DW>++;?=^7>ca+b[
f9Z=\IfVW<_?3Je0WaG[Sd/>ZM]@GK\dDbd^_N.T?4^TYeG,OGSJ-^]X;;(9RU:_
?;:-#V7\R\=.C7Y2YV+>e2F)]#@fbYN,>K0^FW?PNaVE7?+E:M/cPb4a7LJ<<4H7
LReF32^0(I4K?]gdf+HUH9SVCCaMR6C5#T2/KZ8]b.4OS7&\cB_0fY/J/QFFFO#]
bHI1?(ZA]283H&FT8bU.6[EJ24?b5T,=WWSW_f.<g_J]&RQX8Va,5GCF&4T(-X.J
d_c59:9/G\YY<_b-D/Y_]BOZ^(TY^HgA[YCVW9<@WY,dU3QFZ8O6UU;G79CA=_9b
_2OV\&=3+L+Wb.(9KE#4A<QT?eX-CB#=-+CUICgcd:8eJBc(UTG-)Z01(:YEbe(e
X@5HXZUT7E-Ma/1<&0]@aZL[f3QB6?J-Z]LY3W]g)5G_DcIJ6WDAe(L>-K9DaYF[
#Z&+;eHY@[Ud1fWFa:NL?]<YI72f&1NA>g(1SQLJ.+eZ#5:RLBFHG-H/3HIbDQ-A
Z/IHQK,E-C&&G)=^aQ0V3FP9U\CGf\SbMX-I;c43gT?=10YLWF51=2^TWJPO-/P_
4]W>J2.K5<.WGK9SI:93JK6RILQS86+I,T-.JV8IP0:1a:63&?V(@;/R&OMNaE#@
YgbN=BVTXPF:E-_M[O>3NWY1W]\)DV8geDME#1cGJSa6N??,NV>1<Y?^>0V@PbZF
6<BPQT_^+\+&3U5IV-W]C17OEM1/3TJK3(Y6F8/e4YSBTg[-bR6UMZ:4>CDbY?L-
N[gf;PdQH<++ZJbS-KKJ+AV.d1<?;B4;P/V@-LbO0aS7[c&d>=YSVd2EA@IP/J9U
g\HAZLU-+VbL/[F2=Ge@U,d4D^_]MGVO-FN\cYO,-V_&LI[[&eJ?_0eWd2aB[]O2
#W79T5##QGa:P,=Y8JUY^2/.g+NOU&E9-^IKcU:-K--=U:(QZB2T1YWQKdHLM-0_
)+M8fDAIQ_OeMFZ-YaFKQ6a/W.6WU4;eMQbEM/WPC\f>XZNCUe3R82g9<5G_KG0_
48fBINa8Y1JeVL25<KOV>^F;H[?E>ND;@^Y,=@^&0N:\A\ZG2YG#G;eGOG.-7-#F
M#-7F/)[P4:TN9+De)BgI)BG0R-,N(-DI,RU@&@&bEMM^#_JL)WT#1Y[^;190;]d
+<g0I.+,[336]YH-d\Id.]A_[d-]SYYI](.Ic@cNfF)_\Mb>&Y;19#2AUgIKKD(g
I?b+LKUbBG1>1Y?TOdGA@6N#8UBbaRI\g/5=A)\b9/RK]R+J1ZJ-.P\11#T0?T<2
d_GbYEYNTI\;>+;\_EJ;J8>Jg97;Z[/&g;6gPL9\cG#.:0L:I.#I?\f<D&A[eg([
8MSXQ?67YJIgX>;W/W@+[[).M(d]A-(,F\B3K5FRO0@3=g1YS)KLCB(R)VV4?-ZM
,<Z68FMZ1b=&,3Z>9[];d<ME-8K9#Ng1&&aM/;9ZC4=Z66Y10XW=Y?BG1CA_1=ES
-/UP^J<K&7A]fY;K2?g_1S-D]Da=EbG1WQE_9[7e\V8X0>=6?4R..VKFREATGb\K
Xb+d56W(CbN[U1=A?#dPG2:.FHJ?L]N4Pd&cKZgFAQV6bN,bcDWJTW9S;:IR]/BJ
>[dQV?&:ed,Kb(GMV;=KIDfV-@.4KP-(NWO9(f]aZ5gL))3?F[13+R++XQ9APBOY
1W2IQTc9_=O+8A?V.?)4Q^e:_FObL:2c+)G1-MJ-HFCKc/,__]2BUdL)e:LdgdR4
<-@gK.=gF-4bDU3[Q?,IF[F_&_DDLdM8BIV&\7gN3FNS10G+ZRf]eDFWdJBQR8Eg
=1C+[&E=XgYB4A;0#LSZ&?d.DR@(J,-e4gL+58NZVF2N\JW&9K[3\0<(/(aK(8Ce
_#3V0MHb&E[N0;8Tf#HJIgL63FfDbC3fG3M)8AH6#\bU1)7Je/#B]WHc@Yd6<ge)
MY3D+41SJ=:\@T)a3MYQ<GQ:&=&CB/D]W2Ve7+N(DcA<A_+1YFePM-;J7Z]L/:c1
__\=MBBFS\4AD<JAL40J=.PX;9^4MYeQZ(L4/IU1O./U?>CH,XQWaOB0)f:PKOfP
cJcK.[G93YWQB:IHS/-g#b>.FFQ3J(0,D81b_+Tc_=GS&+I/e;(HNJ8g7U9RT5Z.
VQb86LR=Dfc\LX9ddFbZL&2bYJ1\3&W[LY=I1O)[8HA^g7.;D;H\YTc<EBDPB2XR
12:JJ-#>DNZc\OC1^R<gF^D11_,YZI\I^S0fAIIX_]9:6^g9P/Q8(^VD@SE/58]f
Q+dU=_\B8B>e/JAP:LO1P3^C1[bCU@^]Y8\:AZC5V;RBSebbIUe(.:Bb#,P2A0_P
_Ve:#V@P;U0SQ)e;CeAaL(?9d.L<d,50L<LQDgB?DEJ-L.9P><d4=-^C,d@2ab)Y
BKBSI&b^E2d//3:.O77gOH8=&^(aF\BbK@&#()b-T<GGW]3c6IbN;bJ,S6;@F5>C
6PRd7@^^1?GN=[RfP/2QCc<1Gef,,:NZW\+<LG.>Jg:2NBLOFbXaQYeb].91dJR@
HDT51W_AZ)ZCP4Y?USY.YW+9=B<L@<FT?e9O2<2Q>e_g0?ADDf-^:_^V)SE0GKH=
C15^TgDD8+/2LELEa9@-.g3NCSIbX\RXCJ\T\W\4O0dQ=RaIM6@WB1L>JO#T/8FE
##_4J][c?(#I_)8&.]4Z(ZV[Y+<X7dXALFQMbYFL1D+c,UM4R,7P7/Re,e;IC7Jg
>&ff2B-?E7EA8]<+Tc8[D[AO)(;dQCX\,.(2cZX2A?1Y7((DT.W&_VfEWVR9ad1I
1fP;4<_N9DXA,$
`endprotected
endmodule
